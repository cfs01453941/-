# R=RESISTANCE RPERSQ* L/W
RVDD1_1 M6_200000_0  M6_1689000_0 3.7225
RVDD1_2 M6_1689000_0  M6_1689000_359000 0.8975
RVDD1_3 M6_1689000_359000  M6_1698000_359000 0.0225
V_VDD1_1 M6_200000_0 gnd 1
I_VDD1_1 M6_1698000_359000 gnd 0.005

RVDD2_1 M6_19000_500000  M6_1689000_500000 4.175
RVDD2_2 M6_1689000_500000  M6_1689000_549000 0.1225
RVDD2_3 M5_0_500000  M5_19000_500000 0.095
RVDD2_4 M6_1689000_549000  M6_1698000_549000 0.0225
RVDD2_5 M5_19000_500000  M6_19000_500000 5
V_VDD2_1 M5_0_500000 gnd 1
I_VDD2_1 M6_1698000_549000 gnd 0.002

RVDD3_1 M6_0_1019000  M6_1529000_1019000 3.8225
RVDD3_2 M6_1529000_1019000  M6_1529000_1899000 2.2
RVDD3_3 M5_0_1000000  M5_0_1019000 0.095
RVDD3_4 M6_1529000_1899000  M6_1540000_1899000 0.0275
RVDD3_5 M5_0_1019000  M6_0_1019000 5
RVDD3_6 M6_0_991000  M6_0_321000 1.675
RVDD3_7 M6_0_321000  M6_379000_321000 0.9475
RVDD3_8 M5_0_1000000  M5_0_991000 0.045
RVDD3_9 M5_379000_321000  M5_388000_321000 0.045
RVDD3_10 M5_0_991000  M6_0_991000 5
RVDD3_11 M6_379000_321000  M5_379000_321000 5
V_VDD3_1 M5_0_1000000 gnd 1
I_VDD3_1 M6_1540000_1899000 gnd 0.003
I_VDD3_2 M5_388000_321000 gnd 0.002


.tran 1ns 1ns
.end
